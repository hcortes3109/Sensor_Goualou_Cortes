.title KiCad schematic
P1 NC_01 NC_02 NC_03 +3V3 +5V GND GND NC_04 Power
P2 ADC NC_05 NC_06 NC_07 SDA SCK Analog
P5 NC_08 CONN_01X01
P6 NC_09 CONN_01X01
P7 NC_10 CONN_01X01
P8 NC_11 CONN_01X01
P4 NC_12 NC_13 NC_14 CLK DATA SWITCH NC_15 NC_16 Digital
P3 SCK SDA NC_17 GND NC_18 NC_19 TX RX NC_20 NC_21 Digital
R0 +5V Net-_R0-Pad2_ Rsensor
R5 Net-_R0-Pad2_ IN+ 10k
R1 GND IN+ 100k
C1 IN+ GND 100n
R6 ADC Net-_C4-Pad1_ 1k
C2 ADC GND 100n
R2 GND IN- 1k
C4 Net-_C4-Pad1_ IN- 1�
R3 IN- Net-_C4-Pad1_ 100k
C3 +5V GND 100n
U1 NC_22 IN- IN+ GND NC_23 Net-_C4-Pad1_ +5V NC_24 LT1050
U31 +5V GND RX TX Bluetooth-HC05
U41 CLK DATA SWITCH +5V GND KY_040
U21 GND +5V SCK SDA OLED_0.91
.end
